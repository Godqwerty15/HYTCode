module or2(a, b, o);
input a, b;
output o;

assign o = a | b;

endmodule
