module Not2(x, s);
input x;
output s;
assign s = ~x;

endmodule
